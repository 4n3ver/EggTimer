library verilog;
use verilog.vl_types.all;
entity OnBoardTester is
end OnBoardTester;
