library verilog;
use verilog.vl_types.all;
entity ClockDividerTester is
end ClockDividerTester;
